
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY MemIn IS
PORT (
	CLK : IN std_logic; -- clock
	addr : IN integer; -- Address
	WE : IN std_logic; -- Write Enable
	Din : IN integer ; -- Input Data
	RE : IN std_logic; -- Read Enable
	Dout : OUT integer -- Output data
);
END MemIn;

ARCHITECTURE RTL OF MemIn IS
TYPE ARRAY_DATA IS ARRAY (0 TO 1024 - 1) OF Integer;
SIGNAL MemIn_Array : ARRAY_DATA := (
-93, -365, -64, -67, 264, -207, -495, -100, 178, -486, 
-75, -399, 247, -137, 359, 198, 312, -471, -192, 455, -24, 
-492, -283, -29, 136, 199, -12, 1, 350, -66, 19, 210, 495, 
154, -108, -246, 304, 149, 251, -213, -267, 407, -219, -342, 
-264, -159, -305, 304, -176, -201, 440, 389, 474, -100, -469, 
-236, 4, -448, -382, 206, 419, -259, -213, 40, 137, 448, 397, 
321, 86, 131, 46, -309, 487, -81, -3, -2, -89, -225, 50, -443, 
-282, -270, 246, 484, -280, -80, 345, -69, -194, -475, 17, 443, 
43, -80, 411, -16, -205, -75, -418, -429, -326, 76, -230, 352, 
55, -438, -112, -372, 24, 74, 160, -140, -15, 320, -80, 296, 209, 
115, -441, 58, 455, 336, 333, -173, 283, 384, 100, -308, 483, 468, 
177, -379, 84, 286, -164, 468, 43, 270, 454, 27, -135, 463, 365, 138, 
-248, 314, -262, -453, 82, -117, 95, 403, 297, -154, 278, 38, -378, 
359, -86, 191, -60, -296, 275, 421, 138, 181, 58, -66, -70, 170, 73, 
295, 75, 325, -215, -423, 76, 392, 258, 448, 79, -412, -315, -361, 
-40, -461, -261, -161, -337, -277, 121, 274, 214, 328, -20, 186, 
-77, -394, 391, -477, -364, 147, 3, 111, -201, -404, 414, 50, -331, 
226, 382, 417, 356, -180, -35, -268, -419, -434, -442, -169, -288, -5, 
-346, 277, -318, 337, 282, 27, 429, -173, 8, -328, -389, 426, -89, 372, 
-192, -308, -2, 44, -160, -79, 484, -452, 146, 288, -23, 391, -15, 96, 
-236, 342, 290, 28, -219, 259, 395, -432, -387, 420, -448, -320, 294, 
-66, 75, 438, 143, 434, -222, 13, -469, 76, -416, 322, -335, 180, -344, 
426, -491, -217, -280, 263, 290, -188, 155, 16, 153, -482, 199, -330, 319, 
114, -175, -336, -487, 227, -254, -87, -382, -367, -118, -167, -370, 96, 
333, -488, -398, -23, -387, 151, 270, 440, -250, 390, 256, 434, -157, 
-423, -328, 414, 193, -444, -266, -383, 260, -429, -134, 138, -415, 17, 
-366, 142, 464, 16, -484, 86, -441, 133, -375, 274, -439, -25, 263, -472, 
-332, -21, 79, 139, -428, -161, 242, -489, 217, -40, -138, 484, -108, -41, 
-74, -233, -386, -386, 175, -68, -452, 391, -290, 20, -102, 9, -187, 326, 
334, -10, -212, -275, 313, -484, 64, -184, -207, -200, 475, 295, -142, 
175, 431, -302, 341, 56, 116, -352, 395, -206, -390, 178, -331, -333, 
-182, -474, 59, -112, 383, 466, 251, -400, -63, -470, -317, -473, -145, 
147, -286, 84, 464, 171, 83, -379, -125, 350, 351, -385, 31, 187, -412, 
365, -439, -385, -439, 120, -378, -266, -326, 218, -149, 260, -86, -173, 
0, -231, -36, -170, -163, 410, 227, -325, 55, 439, -170, -69, -138, 238, 
-488, 426, -417, 180, -500, 458, -195, -244, 440, -429, 131, 226, -257, 
85, -374, 478, 458, -43, 30, -105, -117, 50, 223, -321, -281, -262, 185, 
-111, -429, -74, -375, -230, -189, 467, -356, 382, -282, 202, 351, 28, 
360, -245, 422, 362, 402, -435, -288, -326, -291, -244, -417, 102, 80, 
-302, 116, 179, 27, 96, 74, -489, -102, 23, -447, 476, -303, -139, -64, 
-213, -14, -213, 228, -212, -209, 406, -61, -393, -382, 492, -348, -28, 
234, -124, 276, -235, -438, 192, -307, 258, -218, -303, -21, 391, -19, 
324, 301, 92, 70, 63, -107, -335, 493, -198, -486, -203, -166, 216, -135, 
480, -2, -71, -201, -360, -391, -460, -453, -333, -16, 340, -400, -255, 
398, 401, 128, 442, -452, -263, -241, -34, -280, 94, 58, 490, 54, 322, 
-215, 119, 289, -108, 460, -377, 211, 355, -62, -498, 436, -145, -382, 
373, -59, -270, -169, 215, -140, -384, -372, -126, -479, 39, 240, 186, 
444, -494, 90, 428, 138, -255, -442, -295, 483, -39, 487, -17, 209, 499, 
39, 171, -441, 218, 331, 174, -344, -316, 326, 15, 460, -86, 108, 466, 
261, -85, 238, 455, -318, 469, 87, -372, -365, 346, 443, 253, -432, -20, 
-462, -51, 402, 55, -356, 165, -371, 379, -10, 134, 210, -481, 271, -453, 
-471, 483, 128, 26, -497, -291, 172, 429, 415, -273, 174, 454, -81, 358, 
-127, -109, -176, -92, 17, -245, 449, 175, -413, 142, -79, 445, 141, 129, 
-7, 279, -35, -170, 228, -192, 305, -171, -418, 365, 56, -160, -20, 369, 56, 
376, -31, -405, -361, 36, 460, 209, 42, 189, -402, -295, -114, 138, 115, 
-476, 135, -111, 265, -417, -347, 91, 289, 317, 488, 417, -267, 64, -371, 
-295, -287, 301, 131, 0, -60, 113, -390, -449, -478, -79, 112, 411, 158, 
-237, 303, -336, -356, -250, 170, -108, 482, 487, -391, 326, -195, 303, 
-160, -103, -94, 23, -492, 95, 288, 205, 87, -265, 463, 44, -322, 341, 
-380, 162, -186, 421, 116, -198, 221, -256, -338, 67, -163, -117, -170, 
447, 21, 490, -97, -78, 166, 181, -497, -453, -385, 298, 114, 97, -148, 
353, -213, -437, -410, 490, -353, 402, 286, 301, -170, 55, -180, 346, 
-472, 74, 275, -277, -195, 425, 324, -134, -318, -231, -290, 109, 285, 
-440, -76, -61, -457, -193, -463, 201, -67, 92, 98, -428, -158, -362, 
433, 116, 352, 380, -177, 188, -471, -498, 21, -299, 392, -54, 462, 33, 
219, -436, 199, -119, 84, 482, -305, 408, 175, 141, 89, -416, -469, -398, 
354, -287, -372, -236, 72, -101, -252, -310, 124, 443, -454, -410, -238, 
-113, 156, 285, 465, -302, 494, 478, -100, -17, 180, 441, -410, -36, -30, 
266, 180, 85, -463, -259, -281, -303, 250, 166, -303, -159, 353, 272, -314, 
-308, -385, 488, -295, -107, 263, 318, 437, 363, 463, -481, -257, 166, -202, 
265, 499, 394, -443, 131, -251, 459, 173, 398, 4, -191, 210, -69, -374, -353, 
35, 226, 162, -468, 483, 417, 205, -213, -291, 313, -376, -52, -14, -446, 225, 
338, 231, 211, 180, -28, 240, 454, -202, -466, -176, -248, -345, -128, -16, 346, 
-232, -3, 32, 295, 240, 325, 136, -73, 499, 308, -66, -31, -241, -300, 92, -474,
18, -447, 260, -52, -57, 231, -314, 135, 447, -341, 387, -3, -291, 394, 469, -195, 
-282, -141, -476, -109, 4, 156, 478, -171, 388, -477, -153, -107, -470, -404, -339, 2, -176, -355
);
BEGIN
-- Read/Write process
RW_Process : PROCESS (CLK)
BEGIN
 IF (CLK'event and CLK = '1') THEN -- rising clock edge
	IF WE = '1' THEN
		MemIn_Array(addr) <= Din;
	ELSIF RE = '1' THEN
		Dout <= MemIn_Array(addr);
	END IF;
 END IF;
END PROCESS RW_Process;
END RTL;